`timescale 1ns / 1ps

module hello_world;
    

initial begin
$display("welcome to verilog");  
$finish;
end


endmodule